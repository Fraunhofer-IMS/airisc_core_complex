../../../airi5c_hasti_constants.vh