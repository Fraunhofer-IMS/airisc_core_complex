//
// Copyright 2022 FRAUNHOFER INSTITUTE OF MICROELECTRONIC CIRCUITS AND SYSTEMS (IMS), DUISBURG, GERMANY.
// --- All rights reserved --- 
// SPDX-License-Identifier: Apache-2.0 WITH SHL-2.1
// Licensed under the Solderpad Hardware License v 2.1 (the “License”);
// you may not use this file except in compliance with the License, or, at your option, the Apache License version 2.0.
// You may obtain a copy of the License at
// https://solderpad.org/licenses/SHL-2.1/
// Unless required by applicable law or agreed to in writing, any work distributed under the License is distributed on an “AS IS” BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and limitations under the License.
//
//
// File              : airi5c_top_asic.v
// Author            : A. Stanitzki
// Creation Date     : 09.10.20
// Version           : 1.0
// Abstract          : AIRI5C top level for the ASIC implementation         
//

`include "airi5c_ctrl_constants.vh"
`include "airi5c_csr_addr_map.vh"
`include "airi5c_hasti_constants.vh"
`include "airi5c_dmi_constants.vh"
`include "airi5c_arch_options.vh"

module airi5c_top_asic(
   input                           clk,
   input                           nreset,
   input                           testmode,
   input                           ext_interrupt,

// scan chain interface for core
/*   input                           sdi,
   output                          sdo,
   input                           sen,*/

// jtag interface
   input                           tdi,
   input                           tck, 
   input                           tms, 
   output                          tdo,

// connections to IMEM/DMEM bus
   output [`HASTI_ADDR_WIDTH-1:0]  imem_haddr,
   output                          imem_hwrite,
   output [`HASTI_SIZE_WIDTH-1:0]  imem_hsize,
   output [`HASTI_BURST_WIDTH-1:0] imem_hburst,
   output                          imem_hmastlock,
   output [`HASTI_PROT_WIDTH-1:0]  imem_hprot,
   output [`HASTI_TRANS_WIDTH-1:0] imem_htrans,
   output [`HASTI_BUS_WIDTH-1:0]   imem_hwdata,
   input  [`HASTI_BUS_WIDTH-1:0]   imem_hrdata,
   input                           imem_hready,
   input                           imem_hresp,
   output [`HASTI_ADDR_WIDTH-1:0]  dmem_haddr,
   output                          dmem_hwrite,
   output [`HASTI_SIZE_WIDTH-1:0]  dmem_hsize,
   output [`HASTI_BURST_WIDTH-1:0] dmem_hburst,
   output                          dmem_hmastlock,
   output [`HASTI_PROT_WIDTH-1:0]  dmem_hprot,
   output [`HASTI_TRANS_WIDTH-1:0] dmem_htrans,
   output [`HASTI_BUS_WIDTH-1:0]   dmem_hwdata,
   input  [`HASTI_BUS_WIDTH-1:0]   dmem_hrdata,
   input                           dmem_hready,
   input                           dmem_hresp,

// -- Chip specific -- 

// GPIOs
   output [7:0]                    oGPIO_D,
   output [7:0]                    oGPIO_EN,
   input  [7:0]                    iGPIO_I,

// UART
   output                          oUART_TX,
   input                           iUART_RX,

// SPI Master
   output                          oSPI1_MOSI,
   input                           iSPI1_MISO,
   output                          oSPI1_SCLK,
   output                          oSPI1_NSS,

// -- Post-Synthesis debug port --
   output reg [7:0]                debug_out
);

  // ndmreset resets everything but the debug module
  wire                            ndmreset;

  // DMI Bus
  // =======
  // signals driven by debug transfer module
  // and received by the debug module  
  wire  [`DMI_ADDR_WIDTH-1:0]     dmi_addr;
  wire  [`DMI_WIDTH-1:0]          dmi_wdata;
  wire  [`DMI_WIDTH-1:0]          dmi_rdata;
  wire                            dmi_en;
  wire                            dmi_wen;
  wire                            dmi_error;
  wire                            dmi_dm_busy;
   
  // Databus- and Peripherybus-Multiplexer signals
  // =============================================
  wire  [`HASTI_BUS_WIDTH-1:0]     muxed_hrdata;
  wire  [`HASTI_RESP_WIDTH-1:0]    muxed_hresp;
  wire                             muxed_hready;
  
  wire [`HASTI_BUS_WIDTH-1:0]     per_hrdata_gpio;
  wire [`HASTI_RESP_WIDTH-1:0]    per_hresp_gpio;
  wire                            per_hready_gpio;
  
  wire [`HASTI_BUS_WIDTH-1:0]     per_hrdata_system_timer;
  wire [`HASTI_RESP_WIDTH-1:0]    per_hresp_system_timer;
  wire                            per_hready_system_timer;
  
  wire [`HASTI_BUS_WIDTH-1:0]     per_hrdata_spi1;
  wire [`HASTI_RESP_WIDTH-1:0]    per_hresp_spi1;
  wire                            per_hready_spi1;
    
  wire [`HASTI_BUS_WIDTH-1:0]     per_hrdata_uart;
  wire [`HASTI_RESP_WIDTH-1:0]    per_hresp_uart;
  wire                            per_hready_uart;    

  wire [`HASTI_BUS_WIDTH-1:0]     per_hrdata_icap;
  wire [`HASTI_RESP_WIDTH-1:0]    per_hresp_icap;
  wire                            per_hready_icap;    
    
  wire                            nrst = nreset & ndmreset;  
  wire                            lock_custom;

  
  // Interrupt signals generated by core local peripherals
  // =====================================================

  wire                            system_timer_tick;

  
  // DMEM bus multiplexer
  // ====================

  airi5c_periph_mux #
  (
    .S_COUNT(6),
    .S_BASE_ADDR({`MEMORY_BASE_ADDR,`SYSTEM_TIMER_BASE_ADDR,`UART1_BASE_ADDR,`SPI1_BASE_ADDR,`GPIO1_BASE_ADDR,`ICAP_BASE_ADDR}),        
    .S_ADDR_WIDTH({`MEMORY_ADDR_WIDTH,`SYSTEM_TIMER_ADDR_WIDTH,`UART1_ADDR_WIDTH,`SPI1_ADDR_WIDTH,`GPIO1_ADDR_WIDTH,`ICAP_ADDR_WIDTH})    
  )
  peripheral_mux ( 
    .clk_i(clk),
    .rst_ni(nrst),
        
    .m_haddr(dmem_haddr),
    .m_hready(muxed_hready),
    .m_hresp(muxed_hresp),
    .m_hrdata(muxed_hrdata), 
    
    .s_hready({dmem_hready,per_hready_system_timer,per_hready_uart,per_hready_spi1,per_hready_gpio,per_hready_icap}),
    .s_hresp({dmem_hresp,per_hresp_system_timer,per_hresp_uart,per_hresp_spi1,per_hresp_gpio,per_hresp_icap}),
    .s_hrdata({dmem_hrdata,per_hrdata_system_timer,per_hrdata_uart,per_hrdata_spi1,per_hrdata_gpio,per_hrdata_icap})
  );

 
  // Core Complex peripherals 
  // ========================

  airi5c_timer #(.BASE_ADDR(`SYSTEM_TIMER_BASE_ADDR)) system_timer
  (
    .nreset(nrst),
    .clk(clk),
  
    .timer_tick(system_timer_tick),

    .haddr(dmem_haddr),
    .hwrite(dmem_hwrite),
    .hsize(dmem_hsize),
    .hburst(dmem_hburst),
    .hmastlock(dmem_hmastlock),
    .hprot(dmem_hprot),
    .htrans(dmem_htrans),
    .hwdata(dmem_hwdata),
    .hrdata(per_hrdata_system_timer),
    .hready(per_hready_system_timer),
    .hresp(per_hresp_system_timer)
  );


  airi5c_gpio #(.BASE_ADDR(`GPIO1_BASE_ADDR),.WIDTH(8)) 
  gpio(
    .nreset(nrst),
    .clk(clk),

    .gpio_d(oGPIO_D),
    .gpio_en(oGPIO_EN),
    .gpio_i(iGPIO_I),

    .haddr(dmem_haddr),
    .hwrite(dmem_hwrite),
    .hsize(dmem_hsize),
    .hburst(dmem_hburst),
    .hmastlock(dmem_hmastlock),
    .hprot(dmem_hprot),
    .htrans(dmem_htrans),
    .hwdata(dmem_hwdata),
    .hrdata(per_hrdata_gpio),
    .hready(per_hready_gpio),
    .hresp(per_hresp_gpio)
  );

  airi5c_uart #(
    .BASE_ADDR(`UART1_BASE_ADDR),
    .TX_ADDR_WIDTH(5),
    .RX_ADDR_WIDTH(5),
    .TX_MARK(8),
    .RX_MARK(24)
  ) uart1
  (
    .n_reset(nrst),
    .clk(clk),

    .tx(oUART_TX), // airi5c to dtm
    .rx(iUART_RX), // dtm to airi5c
    .cts(1'b1),
    .rts(),
  
    .int_any(),
    .int_tx_full(),
    .int_tx_empty(),
    .int_tx_mark_reached(),
    .int_tx_overflow_error(),
    .int_rx_full(),
    .int_rx_empty(),
    .int_rx_mark_reached(),
    .int_rx_overflow_error(),
    .int_rx_underflow_error(),
    .int_rx_noise_error(),
    .int_rx_parity_error(),
    .int_rx_frame_error(),

    .haddr(dmem_haddr),
    .hwrite(dmem_hwrite),
    .htrans(dmem_htrans),
    .hwdata(dmem_hwdata),
    .hrdata(per_hrdata_uart),
    .hready(per_hready_uart),
    .hresp(per_hresp_uart)
  );
  
  airi5c_icap #(
    .BASE_ADDR(`ICAP_BASE_ADDR),
    .CLK_FREQ_HZ(`SYS_CLK_HZ))
  icap1(
    .n_reset(nrst),
    .clk(clk),

    .lock(lock_custom),
    
    .haddr(dmem_haddr),
    .hwrite(dmem_hwrite),
    .hsize(dmem_hsize),
    .hburst(dmem_hburst),
    .hmastlock(dmem_hmastlock),
    .hprot(dmem_hprot),
    .htrans(dmem_htrans),
    .hwdata(dmem_hwdata),
    .hrdata(per_hrdata_icap),
    .hready(per_hready_icap),
    .hresp(per_hresp_icap)
  );
  
  airi5c_spi #(
    .BASE_ADDR(`SPI1_BASE_ADDR),
    .DEFAULT_MASTER(1),
    .DEFAULT_SD(1))
  spi1(
    .n_reset(nrst),
    .clk(clk),
  
    .enable_master(),

    .master_miso(iSPI1_MISO),
    .master_mosi(oSPI1_MOSI),
    .master_sclk(oSPI1_SCLK),
    .master_nss(oSPI1_NSS),

    .slave_miso(),
    .slave_mosi(1'b0),
    .slave_sclk(1'b0),
    .slave_nss(1'b1),

    .haddr(dmem_haddr),
    .hwrite(dmem_hwrite),
    .hsize(dmem_hsize),
    .hburst(dmem_hburst),
    .hmastlock(dmem_hmastlock),
    .hprot(dmem_hprot),
    .htrans(dmem_htrans),
    .hwdata(dmem_hwdata),
    .hrdata(per_hrdata_spi1),
    .hready(per_hready_spi1),
    .hresp(per_hresp_spi1)
  );


// core/hart instances
// ===================
 
airi5c_core airi5c(
  .nreset(nreset),
  .clk(clk),
  .testmode(testmode),

  .ndmreset(ndmreset),
  .ext_interrupts({`N_EXT_INTS{ext_interrupt}}),
  .system_timer_tick(system_timer_tick),
        
  .imem_haddr(imem_haddr),
  .imem_hwrite(imem_hwrite),
  .imem_hsize(imem_hsize),
  .imem_hburst(imem_hburst),
  .imem_hmastlock(imem_hmastlock),
  .imem_hprot(imem_hprot),
  .imem_htrans(imem_htrans),
  .imem_hwdata(imem_hwdata),
  .imem_hrdata(imem_hrdata),
  .imem_hready(imem_hready),
  .imem_hresp(imem_hresp),
         
  .dmem_haddr(dmem_haddr),
  .dmem_hwrite(dmem_hwrite),
  .dmem_hsize(dmem_hsize),
  .dmem_hburst(dmem_hburst),
  .dmem_hmastlock(dmem_hmastlock),
  .dmem_hprot(dmem_hprot),
  .dmem_htrans(dmem_htrans),
  .dmem_hwdata(dmem_hwdata),
  .dmem_hrdata(muxed_hrdata),
  .dmem_hready(muxed_hready), 
  .dmem_hresp(muxed_hresp),
  
  .lock_custom(lock_custom),
  
  .dmi_addr(dmi_addr),
  .dmi_en(dmi_en),
  .dmi_error(dmi_error),
  .dmi_wen(dmi_wen),
  .dmi_wdata(dmi_wdata),
  .dmi_rdata(dmi_rdata),
  .dmi_dm_busy(dmi_dm_busy)
  ); 

// Debug Transfer Module (DTM) 
// ===========================

airi5c_dtm dtm(
  .clk(clk),
  .nreset(nreset),
  .tck(tck),
  .tms(tms),
  .tdi(tdi),
  .tdo(tdo),   
  .dmi_addr(dmi_addr),
  .dmi_en(dmi_en),
  .dmi_error(dmi_error),
  .dmi_wen(dmi_wen),
  .dmi_wdata(dmi_wdata),
  .dmi_rdata(dmi_rdata),
  .dmi_dm_busy(dmi_dm_busy)
);

// Debug port for post-synthesis verification
// ==========================================

reg [31:0] debug_addr;
reg    debug_hwrite;

 // DEBUG Signals
 // =============
 // The debug_out port is used in 
 // verification to output testbench 
 // results from the official ISA tests.
 // It can be handy for silicon verification
 // as well, but might also be excluded from 
 // synthesis.

always @(posedge clk or negedge nreset) begin
  if(~nreset) begin
    debug_out <= 255;
    debug_addr <= 0;
    debug_hwrite <= 1'b0;
  end else begin
    debug_addr <= muxed_hready ? dmem_haddr : debug_addr;
    debug_hwrite <= muxed_hready ? dmem_hwrite : debug_hwrite;
    `ifndef VPIMODE
    if(((debug_addr[7:0] == 8'h00) || (debug_addr == 32'h80010000)) && (debug_hwrite))
    begin
      debug_out <= dmem_hwdata[7:0];
    end
    `endif
    `ifdef VPIMODE
    if((debug_addr == 32'hc0000024) && (debug_hwrite))
    begin     
        //debug_out <= dmem_hwdata[7:0];
        $write("%c",dmem_hwdata[7:0]);
        if((dmem_hwdata[7:0] == 8'h13) || (dmem_hwdata[7:0] == 8'h10)) $fflush(1);
    end
    `endif  
  end
end

endmodule
